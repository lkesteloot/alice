module cyclonev_hps_interface_mpu_general_purpose(
    input wire [31:0] gp_in /* verilator public */,
    output wire [31:0] gp_out /* verilator public */);


endmodule
