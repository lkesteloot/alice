// soc_system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                             //                   clk.clk
		input  wire [28:0] hps_0_f2h_sdram0_data_address,       // hps_0_f2h_sdram0_data.address
		input  wire [7:0]  hps_0_f2h_sdram0_data_burstcount,    //                      .burstcount
		output wire        hps_0_f2h_sdram0_data_waitrequest,   //                      .waitrequest
		output wire [63:0] hps_0_f2h_sdram0_data_readdata,      //                      .readdata
		output wire        hps_0_f2h_sdram0_data_readdatavalid, //                      .readdatavalid
		input  wire        hps_0_f2h_sdram0_data_read,          //                      .read
		input  wire [63:0] hps_0_f2h_sdram0_data_writedata,     //                      .writedata
		input  wire [7:0]  hps_0_f2h_sdram0_data_byteenable,    //                      .byteenable
		input  wire        hps_0_f2h_sdram0_data_write,         //                      .write
		output wire [14:0] memory_mem_a,                        //                memory.mem_a
		output wire [2:0]  memory_mem_ba,                       //                      .mem_ba
		output wire        memory_mem_ck,                       //                      .mem_ck
		output wire        memory_mem_ck_n,                     //                      .mem_ck_n
		output wire        memory_mem_cke,                      //                      .mem_cke
		output wire        memory_mem_cs_n,                     //                      .mem_cs_n
		output wire        memory_mem_ras_n,                    //                      .mem_ras_n
		output wire        memory_mem_cas_n,                    //                      .mem_cas_n
		output wire        memory_mem_we_n,                     //                      .mem_we_n
		output wire        memory_mem_reset_n,                  //                      .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                       //                      .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                      //                      .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                    //                      .mem_dqs_n
		output wire        memory_mem_odt,                      //                      .mem_odt
		output wire [3:0]  memory_mem_dm,                       //                      .mem_dm
		input  wire        memory_oct_rzqin                     //                      .oct_rzqin
	);

	soc_system_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.mem_a                    (memory_mem_a),                        //           memory.mem_a
		.mem_ba                   (memory_mem_ba),                       //                 .mem_ba
		.mem_ck                   (memory_mem_ck),                       //                 .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                     //                 .mem_ck_n
		.mem_cke                  (memory_mem_cke),                      //                 .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                     //                 .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                    //                 .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                    //                 .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                     //                 .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                  //                 .mem_reset_n
		.mem_dq                   (memory_mem_dq),                       //                 .mem_dq
		.mem_dqs                  (memory_mem_dqs),                      //                 .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                    //                 .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                      //                 .mem_odt
		.mem_dm                   (memory_mem_dm),                       //                 .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                    //                 .oct_rzqin
		.h2f_rst_n                (),                                    //        h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                             // f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (hps_0_f2h_sdram0_data_address),       //  f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (hps_0_f2h_sdram0_data_burstcount),    //                 .burstcount
		.f2h_sdram0_WAITREQUEST   (hps_0_f2h_sdram0_data_waitrequest),   //                 .waitrequest
		.f2h_sdram0_READDATA      (hps_0_f2h_sdram0_data_readdata),      //                 .readdata
		.f2h_sdram0_READDATAVALID (hps_0_f2h_sdram0_data_readdatavalid), //                 .readdatavalid
		.f2h_sdram0_READ          (hps_0_f2h_sdram0_data_read),          //                 .read
		.f2h_sdram0_WRITEDATA     (hps_0_f2h_sdram0_data_writedata),     //                 .writedata
		.f2h_sdram0_BYTEENABLE    (hps_0_f2h_sdram0_data_byteenable),    //                 .byteenable
		.f2h_sdram0_WRITE         (hps_0_f2h_sdram0_data_write)          //                 .write
	);

endmodule
